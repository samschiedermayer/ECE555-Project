module mult;

endmodule

