module neuron;

endmodule

