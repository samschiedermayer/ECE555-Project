module adder;

endmodule

